//TODO
module dir_monitor(
  input  wire        clock,
  input  wire[63:0]  id,
  input  wire[7:0]   bus_type,

  input  wire        io_dirWReq_valid,
  input  wire[8:0]   io_dirWReq_bits_set,
  input  wire[2:0]   io_dirWReq_bits_way,
  input  wire        io_dirWReq_bits_data_dirty,
  input  wire[1:0]   io_dirWReq_bits_data_state,
  input  wire[1:0]   io_dirWReq_bits_data_clientStates_0,
  input  wire[1:0]   io_dirWReq_bits_data_clientStates_1,
  input  wire        io_dirWReq_bits_data_prefetch,
  input  wire        io_tagWReq_valid,
  input  wire[8:0]   io_tagWReq_bits_set,
  input  wire[2:0]   io_tagWReq_bits_way,
  input  wire[18:0]  io_tagWReq_bits_tag,
  input  wire        io_clientDirWReq_valid,
  input  wire[6:0]   io_clientDirWReq_bits_set,
  input  wire[2:0]   io_clientDirWReq_bits_way,
  input  wire[1:0]   io_clientDirWReq_bits_data_0_state,
  input  wire[1:0]   io_clientDirWReq_bits_data_0_alias,
  input  wire[1:0]   io_clientDirWReq_bits_data_1_state,
  input  wire[1:0]   io_clientDirWReq_bits_data_1_alias,
  input  wire        io_clientTagWreq_valid,
  input  wire[6:0]   io_clientTagWreq_bits_set,
  input  wire[2:0]   io_clientTagWreq_bits_way,
  input  wire[20:0]  io_clientTagWreq_bits_tag
);

  import "DPI-C" function void dir_monitor_eval(
  input  bit[63:0]  id,
  input  bit[7:0]   bus_type,

  input  bit        io_dirWReq_valid,
  input  bit[8:0]   io_dirWReq_bits_set,
  input  bit[2:0]   io_dirWReq_bits_way,
  input  bit        io_dirWReq_bits_data_dirty,
  input  bit[1:0]   io_dirWReq_bits_data_state,
  input  bit[1:0]   io_dirWReq_bits_data_clientStates_0,
  input  bit[1:0]   io_dirWReq_bits_data_clientStates_1,
  input  bit        io_dirWReq_bits_data_prefetch,
  input  bit        io_tagWReq_valid,
  input  bit[8:0]   io_tagWReq_bits_set,
  input  bit[2:0]   io_tagWReq_bits_way,
  input  bit[18:0]  io_tagWReq_bits_tag,
  input  bit        io_clientDirWReq_valid,
  input  bit[6:0]   io_clientDirWReq_bits_set,
  input  bit[2:0]   io_clientDirWReq_bits_way,
  input  bit[1:0]   io_clientDirWReq_bits_data_0_state,
  input  bit[1:0]   io_clientDirWReq_bits_data_0_alias,
  input  bit[1:0]   io_clientDirWReq_bits_data_1_state,
  input  bit[1:0]   io_clientDirWReq_bits_data_1_alias,
  input  bit        io_clientTagWreq_valid,
  input  bit[6:0]   io_clientTagWreq_bits_set,
  input  bit[2:0]   io_clientTagWreq_bits_way,
  input  bit[20:0]  io_clientTagWreq_bits_tag,
  );

  always@(posedge clock) begin
    dir_monitor_eval(
      id,
      bus_type,

      io_dirWReq_valid,
      io_dirWReq_bits_set,
      io_dirWReq_bits_way,
      io_dirWReq_bits_data_dirty,
      io_dirWReq_bits_data_state,
      io_dirWReq_bits_data_clientStates_0,
      io_dirWReq_bits_data_clientStates_1,
      io_dirWReq_bits_data_prefetch,
      io_tagWReq_valid,
      io_tagWReq_bits_set,
      io_tagWReq_bits_way,
      io_tagWReq_bits_tag,
      io_clientDirWReq_valid,
      io_clientDirWReq_bits_set,
      io_clientDirWReq_bits_way,
      io_clientDirWReq_bits_data_0_state,
      io_clientDirWReq_bits_data_0_alias,
      io_clientDirWReq_bits_data_1_state,
      io_clientDirWReq_bits_data_1_alias,
      io_clientTagWreq_valid,
      io_clientTagWreq_bits_set,
      io_clientTagWreq_bits_way,
      io_clientTagWreq_bits_tag
  );
  end
endmodule